module mem_for_testing(
  input i_clk,
  input [7:0] i_data,
  input [31:0] i_addr,
  input i_write,
  output [7:0] o_data
);

  reg [7:0] memorija[0:511];
  reg [7:0] r_output = 8'd0;

  assign o_data = memorija[i_addr];

  always @(posedge i_clk) begin

    r_output <= memorija[i_addr];
    if (i_write) memorija[i_addr] <= i_data;

  end

  integer i;

  initial begin
   
    for(i = 0; i < 512; i = i + 1)
      memorija[i] = $random;

  end


  wire [7:0] reg0 = memorija[0];
  wire [7:0] reg1 = memorija[1];
  wire [7:0] reg2 = memorija[2];
  wire [7:0] reg3 = memorija[3];
  wire [7:0] reg4 = memorija[4];
  wire [7:0] reg5 = memorija[5];
  wire [7:0] reg6 = memorija[6];
  wire [7:0] reg7 = memorija[7];
  wire [7:0] reg8 = memorija[8];
  wire [7:0] reg9 = memorija[9];
  wire [7:0] reg10 = memorija[10];
  wire [7:0] reg11 = memorija[11];
  wire [7:0] reg12 = memorija[12];
  wire [7:0] reg13 = memorija[13];
  wire [7:0] reg14 = memorija[14];
  wire [7:0] reg15 = memorija[15];
  wire [7:0] reg16 = memorija[16];
  wire [7:0] reg17 = memorija[17];
  wire [7:0] reg18 = memorija[18];
  wire [7:0] reg19 = memorija[19];
  wire [7:0] reg20 = memorija[20];
  wire [7:0] reg21 = memorija[21];
  wire [7:0] reg22 = memorija[22];
  wire [7:0] reg23 = memorija[23];
  wire [7:0] reg24 = memorija[24];
  wire [7:0] reg25 = memorija[25];
  wire [7:0] reg26 = memorija[26];
  wire [7:0] reg27 = memorija[27];
  wire [7:0] reg28 = memorija[28];
  wire [7:0] reg29 = memorija[29];
  wire [7:0] reg30 = memorija[30];
  wire [7:0] reg31 = memorija[31];
  wire [7:0] reg32 = memorija[32];
  wire [7:0] reg33 = memorija[33];
  wire [7:0] reg34 = memorija[34];
  wire [7:0] reg35 = memorija[35];
  wire [7:0] reg36 = memorija[36];
  wire [7:0] reg37 = memorija[37];
  wire [7:0] reg38 = memorija[38];
  wire [7:0] reg39 = memorija[39];
  wire [7:0] reg40 = memorija[40];
  wire [7:0] reg41 = memorija[41];
  wire [7:0] reg42 = memorija[42];
  wire [7:0] reg43 = memorija[43];
  wire [7:0] reg44 = memorija[44];
  wire [7:0] reg45 = memorija[45];
  wire [7:0] reg46 = memorija[46];
  wire [7:0] reg47 = memorija[47];
  wire [7:0] reg48 = memorija[48];
  wire [7:0] reg49 = memorija[49];
  wire [7:0] reg50 = memorija[50];
  wire [7:0] reg51 = memorija[51];
  wire [7:0] reg52 = memorija[52];
  wire [7:0] reg53 = memorija[53];
  wire [7:0] reg54 = memorija[54];
  wire [7:0] reg55 = memorija[55];
  wire [7:0] reg56 = memorija[56];
  wire [7:0] reg57 = memorija[57];
  wire [7:0] reg58 = memorija[58];
  wire [7:0] reg59 = memorija[59];
  wire [7:0] reg60 = memorija[60];
  wire [7:0] reg61 = memorija[61];
  wire [7:0] reg62 = memorija[62];
  wire [7:0] reg63 = memorija[63];
  wire [7:0] reg64 = memorija[64];
  wire [7:0] reg65 = memorija[65];
  wire [7:0] reg66 = memorija[66];
  wire [7:0] reg67 = memorija[67];
  wire [7:0] reg68 = memorija[68];
  wire [7:0] reg69 = memorija[69];
  wire [7:0] reg70 = memorija[70];
  wire [7:0] reg71 = memorija[71];
  wire [7:0] reg72 = memorija[72];
  wire [7:0] reg73 = memorija[73];
  wire [7:0] reg74 = memorija[74];
  wire [7:0] reg75 = memorija[75];
  wire [7:0] reg76 = memorija[76];
  wire [7:0] reg77 = memorija[77];
  wire [7:0] reg78 = memorija[78];
  wire [7:0] reg79 = memorija[79];
  wire [7:0] reg80 = memorija[80];
  wire [7:0] reg81 = memorija[81];
  wire [7:0] reg82 = memorija[82];
  wire [7:0] reg83 = memorija[83];
  wire [7:0] reg84 = memorija[84];
  wire [7:0] reg85 = memorija[85];
  wire [7:0] reg86 = memorija[86];
  wire [7:0] reg87 = memorija[87];
  wire [7:0] reg88 = memorija[88];
  wire [7:0] reg89 = memorija[89];
  wire [7:0] reg90 = memorija[90];
  wire [7:0] reg91 = memorija[91];
  wire [7:0] reg92 = memorija[92];
  wire [7:0] reg93 = memorija[93];
  wire [7:0] reg94 = memorija[94];
  wire [7:0] reg95 = memorija[95];
  wire [7:0] reg96 = memorija[96];
  wire [7:0] reg97 = memorija[97];
  wire [7:0] reg98 = memorija[98];
  wire [7:0] reg99 = memorija[99];
  wire [7:0] reg100 = memorija[100];
  wire [7:0] reg101 = memorija[101];
  wire [7:0] reg102 = memorija[102];
  wire [7:0] reg103 = memorija[103];
  wire [7:0] reg104 = memorija[104];
  wire [7:0] reg105 = memorija[105];
  wire [7:0] reg106 = memorija[106];
  wire [7:0] reg107 = memorija[107];
  wire [7:0] reg108 = memorija[108];
  wire [7:0] reg109 = memorija[109];
  wire [7:0] reg110 = memorija[110];
  wire [7:0] reg111 = memorija[111];
  wire [7:0] reg112 = memorija[112];
  wire [7:0] reg113 = memorija[113];
  wire [7:0] reg114 = memorija[114];
  wire [7:0] reg115 = memorija[115];
  wire [7:0] reg116 = memorija[116];
  wire [7:0] reg117 = memorija[117];
  wire [7:0] reg118 = memorija[118];
  wire [7:0] reg119 = memorija[119];
  wire [7:0] reg120 = memorija[120];
  wire [7:0] reg121 = memorija[121];
  wire [7:0] reg122 = memorija[122];
  wire [7:0] reg123 = memorija[123];
  wire [7:0] reg124 = memorija[124];
  wire [7:0] reg125 = memorija[125];
  wire [7:0] reg126 = memorija[126];
  wire [7:0] reg127 = memorija[127];
  wire [7:0] reg128 = memorija[128];
  wire [7:0] reg129 = memorija[129];
  wire [7:0] reg130 = memorija[130];
  wire [7:0] reg131 = memorija[131];
  wire [7:0] reg132 = memorija[132];
  wire [7:0] reg133 = memorija[133];
  wire [7:0] reg134 = memorija[134];
  wire [7:0] reg135 = memorija[135];
  wire [7:0] reg136 = memorija[136];
  wire [7:0] reg137 = memorija[137];
  wire [7:0] reg138 = memorija[138];
  wire [7:0] reg139 = memorija[139];
  wire [7:0] reg140 = memorija[140];
  wire [7:0] reg141 = memorija[141];
  wire [7:0] reg142 = memorija[142];
  wire [7:0] reg143 = memorija[143];
  wire [7:0] reg144 = memorija[144];
  wire [7:0] reg145 = memorija[145];
  wire [7:0] reg146 = memorija[146];
  wire [7:0] reg147 = memorija[147];
  wire [7:0] reg148 = memorija[148];
  wire [7:0] reg149 = memorija[149];
  wire [7:0] reg150 = memorija[150];
  wire [7:0] reg151 = memorija[151];
  wire [7:0] reg152 = memorija[152];
  wire [7:0] reg153 = memorija[153];
  wire [7:0] reg154 = memorija[154];
  wire [7:0] reg155 = memorija[155];
  wire [7:0] reg156 = memorija[156];
  wire [7:0] reg157 = memorija[157];
  wire [7:0] reg158 = memorija[158];
  wire [7:0] reg159 = memorija[159];
  wire [7:0] reg160 = memorija[160];
  wire [7:0] reg161 = memorija[161];
  wire [7:0] reg162 = memorija[162];
  wire [7:0] reg163 = memorija[163];
  wire [7:0] reg164 = memorija[164];
  wire [7:0] reg165 = memorija[165];
  wire [7:0] reg166 = memorija[166];
  wire [7:0] reg167 = memorija[167];
  wire [7:0] reg168 = memorija[168];
  wire [7:0] reg169 = memorija[169];
  wire [7:0] reg170 = memorija[170];
  wire [7:0] reg171 = memorija[171];
  wire [7:0] reg172 = memorija[172];
  wire [7:0] reg173 = memorija[173];
  wire [7:0] reg174 = memorija[174];
  wire [7:0] reg175 = memorija[175];
  wire [7:0] reg176 = memorija[176];
  wire [7:0] reg177 = memorija[177];
  wire [7:0] reg178 = memorija[178];
  wire [7:0] reg179 = memorija[179];
  wire [7:0] reg180 = memorija[180];
  wire [7:0] reg181 = memorija[181];
  wire [7:0] reg182 = memorija[182];
  wire [7:0] reg183 = memorija[183];
  wire [7:0] reg184 = memorija[184];
  wire [7:0] reg185 = memorija[185];
  wire [7:0] reg186 = memorija[186];
  wire [7:0] reg187 = memorija[187];
  wire [7:0] reg188 = memorija[188];
  wire [7:0] reg189 = memorija[189];
  wire [7:0] reg190 = memorija[190];
  wire [7:0] reg191 = memorija[191];
  wire [7:0] reg192 = memorija[192];
  wire [7:0] reg193 = memorija[193];
  wire [7:0] reg194 = memorija[194];
  wire [7:0] reg195 = memorija[195];
  wire [7:0] reg196 = memorija[196];
  wire [7:0] reg197 = memorija[197];
  wire [7:0] reg198 = memorija[198];
  wire [7:0] reg199 = memorija[199];
  wire [7:0] reg200 = memorija[200];
  wire [7:0] reg201 = memorija[201];
  wire [7:0] reg202 = memorija[202];
  wire [7:0] reg203 = memorija[203];
  wire [7:0] reg204 = memorija[204];
  wire [7:0] reg205 = memorija[205];
  wire [7:0] reg206 = memorija[206];
  wire [7:0] reg207 = memorija[207];
  wire [7:0] reg208 = memorija[208];
  wire [7:0] reg209 = memorija[209];
  wire [7:0] reg210 = memorija[210];
  wire [7:0] reg211 = memorija[211];
  wire [7:0] reg212 = memorija[212];
  wire [7:0] reg213 = memorija[213];
  wire [7:0] reg214 = memorija[214];
  wire [7:0] reg215 = memorija[215];
  wire [7:0] reg216 = memorija[216];
  wire [7:0] reg217 = memorija[217];
  wire [7:0] reg218 = memorija[218];
  wire [7:0] reg219 = memorija[219];
  wire [7:0] reg220 = memorija[220];
  wire [7:0] reg221 = memorija[221];
  wire [7:0] reg222 = memorija[222];
  wire [7:0] reg223 = memorija[223];
  wire [7:0] reg224 = memorija[224];
  wire [7:0] reg225 = memorija[225];
  wire [7:0] reg226 = memorija[226];
  wire [7:0] reg227 = memorija[227];
  wire [7:0] reg228 = memorija[228];
  wire [7:0] reg229 = memorija[229];
  wire [7:0] reg230 = memorija[230];
  wire [7:0] reg231 = memorija[231];
  wire [7:0] reg232 = memorija[232];
  wire [7:0] reg233 = memorija[233];
  wire [7:0] reg234 = memorija[234];
  wire [7:0] reg235 = memorija[235];
  wire [7:0] reg236 = memorija[236];
  wire [7:0] reg237 = memorija[237];
  wire [7:0] reg238 = memorija[238];
  wire [7:0] reg239 = memorija[239];
  wire [7:0] reg240 = memorija[240];
  wire [7:0] reg241 = memorija[241];
  wire [7:0] reg242 = memorija[242];
  wire [7:0] reg243 = memorija[243];
  wire [7:0] reg244 = memorija[244];
  wire [7:0] reg245 = memorija[245];
  wire [7:0] reg246 = memorija[246];
  wire [7:0] reg247 = memorija[247];
  wire [7:0] reg248 = memorija[248];
  wire [7:0] reg249 = memorija[249];
  wire [7:0] reg250 = memorija[250];
  wire [7:0] reg251 = memorija[251];
  wire [7:0] reg252 = memorija[252];
  wire [7:0] reg253 = memorija[253];
  wire [7:0] reg254 = memorija[254];
  wire [7:0] reg255 = memorija[255];
  wire [7:0] reg256 = memorija[256];
  wire [7:0] reg257 = memorija[257];
  wire [7:0] reg258 = memorija[258];
  wire [7:0] reg259 = memorija[259];
  wire [7:0] reg260 = memorija[260];
  wire [7:0] reg261 = memorija[261];
  wire [7:0] reg262 = memorija[262];
  wire [7:0] reg263 = memorija[263];
  wire [7:0] reg264 = memorija[264];
  wire [7:0] reg265 = memorija[265];
  wire [7:0] reg266 = memorija[266];
  wire [7:0] reg267 = memorija[267];
  wire [7:0] reg268 = memorija[268];
  wire [7:0] reg269 = memorija[269];
  wire [7:0] reg270 = memorija[270];
  wire [7:0] reg271 = memorija[271];
  wire [7:0] reg272 = memorija[272];
  wire [7:0] reg273 = memorija[273];
  wire [7:0] reg274 = memorija[274];
  wire [7:0] reg275 = memorija[275];
  wire [7:0] reg276 = memorija[276];
  wire [7:0] reg277 = memorija[277];
  wire [7:0] reg278 = memorija[278];
  wire [7:0] reg279 = memorija[279];
  wire [7:0] reg280 = memorija[280];
  wire [7:0] reg281 = memorija[281];
  wire [7:0] reg282 = memorija[282];
  wire [7:0] reg283 = memorija[283];
  wire [7:0] reg284 = memorija[284];
  wire [7:0] reg285 = memorija[285];
  wire [7:0] reg286 = memorija[286];
  wire [7:0] reg287 = memorija[287];
  wire [7:0] reg288 = memorija[288];
  wire [7:0] reg289 = memorija[289];
  wire [7:0] reg290 = memorija[290];
  wire [7:0] reg291 = memorija[291];
  wire [7:0] reg292 = memorija[292];
  wire [7:0] reg293 = memorija[293];
  wire [7:0] reg294 = memorija[294];
  wire [7:0] reg295 = memorija[295];
  wire [7:0] reg296 = memorija[296];
  wire [7:0] reg297 = memorija[297];
  wire [7:0] reg298 = memorija[298];
  wire [7:0] reg299 = memorija[299];
  wire [7:0] reg300 = memorija[300];
  wire [7:0] reg301 = memorija[301];
  wire [7:0] reg302 = memorija[302];
  wire [7:0] reg303 = memorija[303];
  wire [7:0] reg304 = memorija[304];
  wire [7:0] reg305 = memorija[305];
  wire [7:0] reg306 = memorija[306];
  wire [7:0] reg307 = memorija[307];
  wire [7:0] reg308 = memorija[308];
  wire [7:0] reg309 = memorija[309];
  wire [7:0] reg310 = memorija[310];
  wire [7:0] reg311 = memorija[311];
  wire [7:0] reg312 = memorija[312];
  wire [7:0] reg313 = memorija[313];
  wire [7:0] reg314 = memorija[314];
  wire [7:0] reg315 = memorija[315];
  wire [7:0] reg316 = memorija[316];
  wire [7:0] reg317 = memorija[317];
  wire [7:0] reg318 = memorija[318];
  wire [7:0] reg319 = memorija[319];
  wire [7:0] reg320 = memorija[320];
  wire [7:0] reg321 = memorija[321];
  wire [7:0] reg322 = memorija[322];
  wire [7:0] reg323 = memorija[323];
  wire [7:0] reg324 = memorija[324];
  wire [7:0] reg325 = memorija[325];
  wire [7:0] reg326 = memorija[326];
  wire [7:0] reg327 = memorija[327];
  wire [7:0] reg328 = memorija[328];
  wire [7:0] reg329 = memorija[329];
  wire [7:0] reg330 = memorija[330];
  wire [7:0] reg331 = memorija[331];
  wire [7:0] reg332 = memorija[332];
  wire [7:0] reg333 = memorija[333];
  wire [7:0] reg334 = memorija[334];
  wire [7:0] reg335 = memorija[335];
  wire [7:0] reg336 = memorija[336];
  wire [7:0] reg337 = memorija[337];
  wire [7:0] reg338 = memorija[338];
  wire [7:0] reg339 = memorija[339];
  wire [7:0] reg340 = memorija[340];
  wire [7:0] reg341 = memorija[341];
  wire [7:0] reg342 = memorija[342];
  wire [7:0] reg343 = memorija[343];
  wire [7:0] reg344 = memorija[344];
  wire [7:0] reg345 = memorija[345];
  wire [7:0] reg346 = memorija[346];
  wire [7:0] reg347 = memorija[347];
  wire [7:0] reg348 = memorija[348];
  wire [7:0] reg349 = memorija[349];
  wire [7:0] reg350 = memorija[350];
  wire [7:0] reg351 = memorija[351];
  wire [7:0] reg352 = memorija[352];
  wire [7:0] reg353 = memorija[353];
  wire [7:0] reg354 = memorija[354];
  wire [7:0] reg355 = memorija[355];
  wire [7:0] reg356 = memorija[356];
  wire [7:0] reg357 = memorija[357];
  wire [7:0] reg358 = memorija[358];
  wire [7:0] reg359 = memorija[359];
  wire [7:0] reg360 = memorija[360];
  wire [7:0] reg361 = memorija[361];
  wire [7:0] reg362 = memorija[362];
  wire [7:0] reg363 = memorija[363];
  wire [7:0] reg364 = memorija[364];
  wire [7:0] reg365 = memorija[365];
  wire [7:0] reg366 = memorija[366];
  wire [7:0] reg367 = memorija[367];
  wire [7:0] reg368 = memorija[368];
  wire [7:0] reg369 = memorija[369];
  wire [7:0] reg370 = memorija[370];
  wire [7:0] reg371 = memorija[371];
  wire [7:0] reg372 = memorija[372];
  wire [7:0] reg373 = memorija[373];
  wire [7:0] reg374 = memorija[374];
  wire [7:0] reg375 = memorija[375];
  wire [7:0] reg376 = memorija[376];
  wire [7:0] reg377 = memorija[377];
  wire [7:0] reg378 = memorija[378];
  wire [7:0] reg379 = memorija[379];
  wire [7:0] reg380 = memorija[380];
  wire [7:0] reg381 = memorija[381];
  wire [7:0] reg382 = memorija[382];
  wire [7:0] reg383 = memorija[383];
  wire [7:0] reg384 = memorija[384];
  wire [7:0] reg385 = memorija[385];
  wire [7:0] reg386 = memorija[386];
  wire [7:0] reg387 = memorija[387];
  wire [7:0] reg388 = memorija[388];
  wire [7:0] reg389 = memorija[389];
  wire [7:0] reg390 = memorija[390];
  wire [7:0] reg391 = memorija[391];
  wire [7:0] reg392 = memorija[392];
  wire [7:0] reg393 = memorija[393];
  wire [7:0] reg394 = memorija[394];
  wire [7:0] reg395 = memorija[395];
  wire [7:0] reg396 = memorija[396];
  wire [7:0] reg397 = memorija[397];
  wire [7:0] reg398 = memorija[398];
  wire [7:0] reg399 = memorija[399];
  wire [7:0] reg400 = memorija[400];
  wire [7:0] reg401 = memorija[401];
  wire [7:0] reg402 = memorija[402];
  wire [7:0] reg403 = memorija[403];
  wire [7:0] reg404 = memorija[404];
  wire [7:0] reg405 = memorija[405];
  wire [7:0] reg406 = memorija[406];
  wire [7:0] reg407 = memorija[407];
  wire [7:0] reg408 = memorija[408];
  wire [7:0] reg409 = memorija[409];
  wire [7:0] reg410 = memorija[410];
  wire [7:0] reg411 = memorija[411];
  wire [7:0] reg412 = memorija[412];
  wire [7:0] reg413 = memorija[413];
  wire [7:0] reg414 = memorija[414];
  wire [7:0] reg415 = memorija[415];
  wire [7:0] reg416 = memorija[416];
  wire [7:0] reg417 = memorija[417];
  wire [7:0] reg418 = memorija[418];
  wire [7:0] reg419 = memorija[419];
  wire [7:0] reg420 = memorija[420];
  wire [7:0] reg421 = memorija[421];
  wire [7:0] reg422 = memorija[422];
  wire [7:0] reg423 = memorija[423];
  wire [7:0] reg424 = memorija[424];
  wire [7:0] reg425 = memorija[425];
  wire [7:0] reg426 = memorija[426];
  wire [7:0] reg427 = memorija[427];
  wire [7:0] reg428 = memorija[428];
  wire [7:0] reg429 = memorija[429];
  wire [7:0] reg430 = memorija[430];
  wire [7:0] reg431 = memorija[431];
  wire [7:0] reg432 = memorija[432];
  wire [7:0] reg433 = memorija[433];
  wire [7:0] reg434 = memorija[434];
  wire [7:0] reg435 = memorija[435];
  wire [7:0] reg436 = memorija[436];
  wire [7:0] reg437 = memorija[437];
  wire [7:0] reg438 = memorija[438];
  wire [7:0] reg439 = memorija[439];
  wire [7:0] reg440 = memorija[440];
  wire [7:0] reg441 = memorija[441];
  wire [7:0] reg442 = memorija[442];
  wire [7:0] reg443 = memorija[443];
  wire [7:0] reg444 = memorija[444];
  wire [7:0] reg445 = memorija[445];
  wire [7:0] reg446 = memorija[446];
  wire [7:0] reg447 = memorija[447];
  wire [7:0] reg448 = memorija[448];
  wire [7:0] reg449 = memorija[449];
  wire [7:0] reg450 = memorija[450];
  wire [7:0] reg451 = memorija[451];
  wire [7:0] reg452 = memorija[452];
  wire [7:0] reg453 = memorija[453];
  wire [7:0] reg454 = memorija[454];
  wire [7:0] reg455 = memorija[455];
  wire [7:0] reg456 = memorija[456];
  wire [7:0] reg457 = memorija[457];
  wire [7:0] reg458 = memorija[458];
  wire [7:0] reg459 = memorija[459];
  wire [7:0] reg460 = memorija[460];
  wire [7:0] reg461 = memorija[461];
  wire [7:0] reg462 = memorija[462];
  wire [7:0] reg463 = memorija[463];
  wire [7:0] reg464 = memorija[464];
  wire [7:0] reg465 = memorija[465];
  wire [7:0] reg466 = memorija[466];
  wire [7:0] reg467 = memorija[467];
  wire [7:0] reg468 = memorija[468];
  wire [7:0] reg469 = memorija[469];
  wire [7:0] reg470 = memorija[470];
  wire [7:0] reg471 = memorija[471];
  wire [7:0] reg472 = memorija[472];
  wire [7:0] reg473 = memorija[473];
  wire [7:0] reg474 = memorija[474];
  wire [7:0] reg475 = memorija[475];
  wire [7:0] reg476 = memorija[476];
  wire [7:0] reg477 = memorija[477];
  wire [7:0] reg478 = memorija[478];
  wire [7:0] reg479 = memorija[479];
  wire [7:0] reg480 = memorija[480];
  wire [7:0] reg481 = memorija[481];
  wire [7:0] reg482 = memorija[482];
  wire [7:0] reg483 = memorija[483];
  wire [7:0] reg484 = memorija[484];
  wire [7:0] reg485 = memorija[485];
  wire [7:0] reg486 = memorija[486];
  wire [7:0] reg487 = memorija[487];
  wire [7:0] reg488 = memorija[488];
  wire [7:0] reg489 = memorija[489];
  wire [7:0] reg490 = memorija[490];
  wire [7:0] reg491 = memorija[491];
  wire [7:0] reg492 = memorija[492];
  wire [7:0] reg493 = memorija[493];
  wire [7:0] reg494 = memorija[494];
  wire [7:0] reg495 = memorija[495];
  wire [7:0] reg496 = memorija[496];
  wire [7:0] reg497 = memorija[497];
  wire [7:0] reg498 = memorija[498];
  wire [7:0] reg499 = memorija[499];
  wire [7:0] reg500 = memorija[500];
  wire [7:0] reg501 = memorija[501];
  wire [7:0] reg502 = memorija[502];
  wire [7:0] reg503 = memorija[503];
  wire [7:0] reg504 = memorija[504];
  wire [7:0] reg505 = memorija[505];
  wire [7:0] reg506 = memorija[506];
  wire [7:0] reg507 = memorija[507];
  wire [7:0] reg508 = memorija[508];
  wire [7:0] reg509 = memorija[509];
  wire [7:0] reg510 = memorija[510];
  wire [7:0] reg511 = memorija[511];

endmodule
